//=========================================================
// RISC-V SINGLE-CYCLE PROCESSOR
//=========================================================
//
// - Implements basic RV32I subset (User ISA v2.2, May 2017)
// - Supports load/store, R-type, I-type, branch, and jump
// - Extended with custom instructions (ANDN, ORN, XNOR, MIN, MAX, etc.)
// - Designed for simulation using testbench below
// - "Simulation succeeded" when memory[100] = 25
//
//=========================================================
// Author: Sanket Daduria
//=========================================================

module testbench();

  logic clk;
  logic reset;

  logic [31:0] WriteData, DataAdr;
  logic MemWrite;

  // Instantiate the top-level processor system
  top dut(clk, reset, WriteData, DataAdr, MemWrite);
  
  // Initialize reset
  initial begin
    reset <= 1; #22; reset <= 0;
  end

  // Generate waveform for debugging
  initial begin
    $dumpfile("wave.vcd");
    $dumpvars(0, testbench);
  end

  // Clock generation (10ns period)
  always begin
    clk <= 1; #5; clk <= 0; #5;
  end

  // Monitor memory writes to verify simulation result
  always @(negedge clk) begin
    if (MemWrite) begin
      if (DataAdr === 100 && WriteData === 25) begin
        $display("Simulation succeeded");
        $stop;
      end else if (DataAdr !== 96) begin
        $display("Simulation failed");
        $stop;
      end
    end
  end
endmodule


//=========================================================
// TOP MODULE: connects processor core with instruction/data memory
//=========================================================
module top(input  logic clk, reset, 
           output logic [31:0] WriteData, DataAdr, 
           output logic MemWrite);

  logic [31:0] PC, Instr, ReadData;
  
  // Instantiate core and memories
  riscvsingle rvsingle(clk, reset, PC, Instr, MemWrite, DataAdr, 
                       WriteData, ReadData);
  imem imem(PC, Instr);
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);
endmodule


//=========================================================
// RISC-V SINGLE-CYCLE CPU
//=========================================================
module riscvsingle(input  logic clk, reset,
                   output logic [31:0] PC,
                   input  logic [31:0] Instr,
                   output logic MemWrite,
                   output logic [31:0] ALUResult, WriteData,
                   input  logic [31:0] ReadData);

  logic ALUSrc, RegWrite, Jump, Zero;
  logic [1:0] ResultSrc, ImmSrc;
  logic [3:0] ALUControl;

  // Controller generates control signals
  controller c(Instr[6:0], Instr[14:12], Instr[30], Instr[26:25], Zero,
               ResultSrc, MemWrite, PCSrc,
               ALUSrc, RegWrite, Jump,
               ImmSrc, ALUControl);

  // Datapath performs data operations
  datapath dp(clk, reset, ResultSrc, PCSrc,
              ALUSrc, RegWrite,
              ImmSrc, ALUControl,
              Zero, PC, Instr,
              ALUResult, WriteData, ReadData);
endmodule


//=========================================================
// CONTROLLER: Generates control signals for datapath
//=========================================================
module controller(input  logic [6:0] op,
                  input  logic [2:0] funct3,
                  input  logic       funct7b5,
                  input  logic [1:0] funct7b10, 
                  input  logic       Zero,
                  output logic [1:0] ResultSrc,
                  output logic       MemWrite,
                  output logic       PCSrc, ALUSrc,
                  output logic       RegWrite, Jump,
                  output logic [1:0] ImmSrc,
                  output logic [3:0] ALUControl);

  logic [1:0] ALUOp;
  logic Branch;

  // Main decoder: instruction type decoding
  maindec md(op, ResultSrc, MemWrite, Branch,
             ALUSrc, RegWrite, Jump, ImmSrc, ALUOp);

  // ALU decoder: selects ALU operation based on funct fields
  aludec  ad(op[5], funct3, funct7b5, funct7b10, ALUOp, ALUControl);

  // Program Counter select logic
  assign PCSrc = (Branch & Zero) | Jump;
endmodule


//=========================================================
// MAIN DECODER: Decodes opcode to control signals
//=========================================================
module maindec(input  logic [6:0] op,
               output logic [1:0] ResultSrc,
               output logic       MemWrite,
               output logic       Branch, ALUSrc,
               output logic       RegWrite, Jump,
               output logic [1:0] ImmSrc,
               output logic [1:0] ALUOp);

  logic [10:0] controls;

  assign {RegWrite, ImmSrc, ALUSrc, MemWrite,
          ResultSrc, Branch, ALUOp, Jump} = controls;

  always_comb
    case(op)
      //            RW  IS AL MW RS BR AO J
      7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
      7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
      7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type
      7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
      7'b0010011: controls = 11'b1_00_1_0_00_0_10_0; // I-type ALU
      7'b1101111: controls = 11'b1_11_0_0_10_0_00_1; // jal
      7'b0001011: controls = 11'b1_xx_0_0_00_0_11_0; // custom R-type (new ops)
      default:    controls = 11'bx_xx_x_x_xx_x_xx_x; // undefined instruction
    endcase
endmodule


//=========================================================
// ALU DECODER: Determines ALUControl signal
//=========================================================
module aludec(input  logic       opb5,
              input  logic [2:0] funct3,
              input  logic       funct7b5, 
              input  logic [1:0] funct7b10, 
              input  logic [1:0] ALUOp,
              output logic [3:0] ALUControl);

  logic RtypeSub;
  assign RtypeSub = funct7b5 & opb5; // identifies SUB instruction

  always_comb
    case(ALUOp)
      2'b00: ALUControl = 4'b0000; // addition
      2'b01: ALUControl = 4'b0001; // subtraction
      2'b10: case(funct3)
               3'b000: ALUControl = RtypeSub ? 4'b0001 : 4'b0000; // add/sub
               3'b010: ALUControl = 4'b0101; // slt/slti
               3'b110: ALUControl = 4'b0011; // or/ori
               3'b111: ALUControl = 4'b0010; // and/andi
               default: ALUControl = 4'bxxxx;
             endcase
      default: case({funct7b10,funct3})
                 {2'b00, 3'b000}: ALUControl = 4'b0110; // ANDN
                 {2'b00, 3'b001}: ALUControl = 4'b0111; // ORN
                 {2'b00, 3'b010}: ALUControl = 4'b1000; // XNOR
                 {2'b01, 3'b000}: ALUControl = 4'b1001; // MIN
                 {2'b01, 3'b001}: ALUControl = 4'b1010; // MAX
                 {2'b01, 3'b010}: ALUControl = 4'b1011; // MINU
                 {2'b01, 3'b011}: ALUControl = 4'b1100; // MAXU
                 {2'b10, 3'b000}: ALUControl = 4'b1101; // ROL
                 {2'b10, 3'b001}: ALUControl = 4'b1110; // ROR
                 {2'b11, 3'b000}: ALUControl = 4'b1111; // ABS
                 default:          ALUControl = 4'bxxxx;
               endcase
    endcase
endmodule


//=========================================================
// DATAPATH: Connects registers, ALU, PC, and memory
//=========================================================
module datapath(input  logic clk, reset,
                input  logic [1:0]  ResultSrc, 
                input  logic        PCSrc, ALUSrc,
                input  logic        RegWrite,
                input  logic [1:0]  ImmSrc,
                input  logic [3:0]  ALUControl,
                output logic        Zero,
                output logic [31:0] PC,
                input  logic [31:0] Instr,
                output logic [31:0] ALUResult, WriteData,
                input  logic [31:0] ReadData);

  logic [31:0] PCNext, PCPlus4, PCTarget;
  logic [31:0] ImmExt;
  logic [31:0] SrcA, SrcB;
  logic [31:0] Result;

  // Next PC logic
  flopr #(32) pcreg(clk, reset, PCNext, PC); 
  adder       pcadd4(PC, 32'd4, PCPlus4);
  adder       pcaddbranch(PC, ImmExt, PCTarget);
  mux2 #(32)  pcmux(PCPlus4, PCTarget, PCSrc, PCNext);
 
  // Register file read/write
  regfile     rf(clk, RegWrite, Instr[19:15], Instr[24:20], 
                 Instr[11:7], Result, SrcA, WriteData);

  // Immediate generation
  extend      ext(Instr[31:7], ImmSrc, ImmExt);

  // ALU operation
  mux2 #(32)  srcbmux(WriteData, ImmExt, ALUSrc, SrcB);
  alu         alu(SrcA, SrcB, ALUControl, ALUResult, Zero);

  // Result selection: ALU result / memory data / PC+4
  mux3 #(32)  resultmux(ALUResult, ReadData, PCPlus4, ResultSrc, Result);
endmodule


//=========================================================
// REGISTER FILE
//=========================================================
module regfile(input  logic clk, 
               input  logic we3, 
               input  logic [4:0] a1, a2, a3, 
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0]; // 32 registers

  // Write on rising edge if write enabled and not x0
  always_ff @(posedge clk)
    if (we3 & (a3 != 0)) rf[a3] <= wd3;

  // Read ports are combinational
  assign rd1 = (a1 != 0) ? rf[a1] : 0;
  assign rd2 = (a2 != 0) ? rf[a2] : 0;
endmodule


//=========================================================
// SIMPLE ADDER
//=========================================================
module adder(input  [31:0] a, b,
             output [31:0] y);
  assign y = a + b;
endmodule


//=========================================================
// IMMEDIATE EXTENSION UNIT
//=========================================================
module extend(input  logic [31:7] instr,
              input  logic [1:0]  immsrc,
              output logic [31:0] immext);
 
  always_comb
    case(immsrc)
      2'b00: immext = {{20{instr[31]}}, instr[31:20]};              // I-type
      2'b01: immext = {{20{instr[31]}}, instr[31:25], instr[11:7]}; // S-type
      2'b10: immext = {{20{instr[31]}}, instr[7], instr[30:25],
                        instr[11:8], 1'b0};                         // B-type
      2'b11: immext = {{12{instr[31]}}, instr[19:12], instr[20],
                        instr[30:21], 1'b0};                        // J-type
      default: immext = 32'bx;
    endcase             
endmodule


//=========================================================
// GENERIC REGISTER (FLIP-FLOP WITH RESET)
//=========================================================
module flopr #(parameter WIDTH = 8)
              (input  logic clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule


//=========================================================
// MUXES
//=========================================================
module mux2 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, 
              input  logic s, 
              output logic [WIDTH-1:0] y);
  assign y = s ? d1 : d0; 
endmodule

module mux3 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, d2,
              input  logic [1:0] s, 
              output logic [WIDTH-1:0] y);
  assign y = s[1] ? d2 : (s[0] ? d1 : d0); 
endmodule


//=========================================================
// INSTRUCTION MEMORY (read-only, preloaded from riscvtest.hex)
//=========================================================
module imem(input  logic [31:0] a,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0];

  initial $readmemh("riscvtest.hex", RAM);

  assign rd = RAM[a[31:2]]; // word-aligned access
endmodule


//=========================================================
// DATA MEMORY (word-aligned read/write)
//=========================================================
module dmem(input  logic clk, we,
            input  logic [31:0] a, wd,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0];

  assign rd = RAM[a[31:2]];

  always_ff @(posedge clk)
    if (we) RAM[a[31:2]] <= wd;
endmodule


//=========================================================
// ALU: Performs arithmetic, logic, and custom ops
//=========================================================
module alu(input  logic [31:0] a, b,
           input  logic [3:0]  alucontrol,
           output logic [31:0] result,
           output logic        zero);

  logic [31:0] condinvb, sum;
  logic v;              // overflow
  logic isAddSub;       // flag for add/sub
  logic [4:0] shamt;    // shift amount for ROL/ROR

  // Prepare operands for add/sub
  assign condinvb = alucontrol[0] ? ~b : b;
  assign sum = a + condinvb + alucontrol[0];
  assign isAddSub = ~alucontrol[2] & ~alucontrol[1] |
                    ~alucontrol[1] & alucontrol[0];
  assign shamt = b[4:0];

  always_comb
    case (alucontrol)
      4'b0000: result = sum;                                  // ADD
      4'b0001: result = sum;                                  // SUB  
      4'b0010: result = a & b;                                // AND
      4'b0011: result = a | b;                                // OR 
      4'b0100: result = a ^ b;                                // XOR
      4'b0101: result = sum[31] ^ v;                          // SLT
      4'b0110: result = (a & (~b));                           // ANDN
      4'b0111: result = (a | (~b));                           // ORN
      4'b1000: result = ~(a ^ b);                             // XNOR 
      4'b1001: result = (($signed(a) < $signed(b)) ? a : b);  // MIN
      4'b1010: result = (($signed(a) > $signed(b)) ? a : b);  // MAX
      4'b1011: result = ((a < b) ? a : b);                    // MINU
      4'b1100: result = ((a > b) ? a : b);                    // MAXU
      4'b1101: result = (a << shamt) | (a >> (32 - shamt));   // ROL
      4'b1110: result = (a >> shamt) | (a << (32 - shamt));   // ROR
      4'b1111: result = (a[31] == 1'b0) ? a : -a;             // ABS
      default: result = 32'bx;
    endcase

  assign zero = (result == 32'b0);
  assign v = ~(alucontrol[0] ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;
  
endmodule



// Single-cycle implementation of RISC-V (RV32I)
// User-level Instruction Set Architecture V2.2 (May 7, 2017)
// Implements a subset of the base integer instructions:
//    lw, sw
//    add, sub, and, or, slt, 
//    addi, andi, ori, slti
//    beq
//    jal
// Exceptions, traps, and interrupts not implemented
// little-endian memory

// 31 32-bit registers x1-x31, x0 hardwired to 0
// R-Type instructions
//   add, sub, and, or, slt
//   INSTR rd, rs1, rs2
//   Instr[31:25] = funct7 (funct7b5 & opb5 = 1 for sub, 0 for others)
//   Instr[24:20] = rs2
//   Instr[19:15] = rs1
//   Instr[14:12] = funct3
//   Instr[11:7]  = rd
//   Instr[6:0]   = opcode
// I-Type Instructions
//   lw, I-type ALU (addi, andi, ori, slti)
//   lw:         INSTR rd, imm(rs1)
//   I-type ALU: INSTR rd, rs1, imm (12-bit signed)
//   Instr[31:20] = imm[11:0]
//   Instr[24:20] = rs2
//   Instr[19:15] = rs1
//   Instr[14:12] = funct3
//   Instr[11:7]  = rd
//   Instr[6:0]   = opcode
// S-Type Instruction
//   sw rs2, imm(rs1) (store rs2 into address specified by rs1 + immm)
//   Instr[31:25] = imm[11:5] (offset[11:5])
//   Instr[24:20] = rs2 (src)
//   Instr[19:15] = rs1 (base)
//   Instr[14:12] = funct3
//   Instr[11:7]  = imm[4:0]  (offset[4:0])
//   Instr[6:0]   = opcode
// B-Type Instruction
//   beq rs1, rs2, imm (PCTarget = PC + (signed imm x 2))
//   Instr[31:25] = imm[12], imm[10:5]
//   Instr[24:20] = rs2
//   Instr[19:15] = rs1
//   Instr[14:12] = funct3
//   Instr[11:7]  = imm[4:1], imm[11]
//   Instr[6:0]   = opcode
// J-Type Instruction
//   jal rd, imm  (signed imm is multiplied by 2 and added to PC, rd = PC+4)
//   Instr[31:12] = imm[20], imm[10:1], imm[11], imm[19:12]
//   Instr[11:7]  = rd
//   Instr[6:0]   = opcode

//   Instruction  opcode    funct3    funct7
//   sub          0110011   000       0100000
//   add          0110011   000       0000000
//   addi         0010011   000       immediate
//   and          0110011   111       0000000
//   andi         0010011   111       immediate
//   or           0110011   110       000000
//   ori          0010011   110       immediate
//   slt          0110011   010       0000000
//   slti         0010011   010       immediate
//   beq          1100011   000       immediate
//   lw	          0000011   010       immediate
//   sw           0100011   010       immediate
//   jal          1101111   immediate immediate
